��k-      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby��wzrost�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��h2�f8�����R�(KhHNNNJ����J����K t�b�C              �?�t�bhLh&�scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hK�
node_count�K	�nodes�h(h+K ��h-��R�(KK	��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hxhGK ��hyhGK��hzhGK��h{hXK��h|hXK ��h}hGK(��h~hXK0��uK8KKt�b�B�                              @     ��?             H@������������������������       �                     9@                          �E@���}<S�?             7@                            @z�G�z�?	             $@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@�t�b�values�h(h+K ��h-��R�(KK	KK��hX�C�      ;@      5@      9@               @      5@       @       @       @      �?              �?       @                      @              *@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                              @�q�q��?!             H@������������������������       �        	             ,@       
                     @��hJ,�?             A@       	                    @�eP*L��?	             &@                          �@@r�q��?             @������������������������       �                     @                           C@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     7@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      3@      =@      ,@              @      =@      @      @      @      �?      @               @      �?              �?       @                      @              7@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @�q�q��?             H@������������������������       �                     .@                            @<���D�?            �@@                          Pf@X�<ݚ�?             "@������������������������       �                     @                           C@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      3@      =@      .@              @      =@      @      @              @      @       @               @      @                      8@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @�q���?             H@������������������������       �                     3@                            @\-��p�?             =@                        �<eZ@�q�q�?             (@������������������������       �                      @                           h@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     1@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      7@      9@      3@              @      9@      @       @       @               @       @               @       @                      1@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @�q�q�?#             H@������������������������       �                     2@                            @��S�ۿ?             >@                          �0@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      4@      <@      2@               @      <@       @      @       @                      @              8@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                             '@     ��?             H@������������������������       �                      @                           @(옄��?             G@                            @�4�����?             ?@       
                    C@���7�?             6@                            @�����H�?             "@������������������������       �                     @       	                   �@@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             *@������������������������       �                     "@������������������������       �                     .@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      5@      ;@               @      5@      9@      5@      $@      5@      �?       @      �?      @              @      �?      @                      �?      *@                      "@              .@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                            �e@�q�q�?             H@                            @�q�q�?             "@������������������������       �                     @������������������������       �                     @                            @��Sݭg�?            �C@                           @�q�q�?	             .@       
                   �g@�C��2(�?             &@       	                    C@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     8@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      0@      @@      @      @      @                      @      $@      =@      $@      @      $@      �?       @      �?              �?       @               @                      @              8@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @      �?             H@������������������������       �                     4@                          @@@؇���X�?             <@                            @      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     4@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      8@      8@      4@              @      8@      @      @      @                      @              4@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�         
                  y
F@r�qG�?             H@                            @     ��?             @@������������������������       �                     @       	                     @ ��WV�?             :@                           @r�q��?             @                          �0@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     4@                           �?      �?
             0@������������������������       �                     $@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      1@      ?@      @      9@      @              �?      9@      �?      @      �?       @      �?                       @              @              4@      $@      @      $@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                              @r�q��?             H@������������������������       �        
             3@                          �0@ܷ��?��?             =@                           '@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �h@ ��WV�?             :@������������������������       �                     3@	       
                     @؇���X�?             @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      6@      :@      3@              @      :@       @      �?              �?       @              �?      9@              3@      �?      @      �?                      @�t�bubhhubehhub.